red <= NOT ball_on(0) AND NOT ball_on(3) AND NOT ball_on(6) AND NOT ball_on(9) AND NOT cursor_on NOT ball_on(12) AND NOT ball_on(15) AND NOT ball_on(18) AND NOT ball_on(21) AND NOT ball_on(24) AND NOT ball_on(27) AND NOT ball_on(30) AND NOT ball_on(33) AND NOT ball_on(36) AND NOT ball_on(39) AND NOT ball_on(42) AND NOT ball_on(45);
    blue <= NOT ball_on(1) AND NOT ball_on(4) AND NOT ball_on(7) AND NOT ball_on(10) AND NOT cursor_on NOT ball_on(13) AND NOT ball_on(16) AND NOT ball_on(19) AND NOT ball_on(22) AND NOT ball_on(25) AND NOT ball_on(28) AND NOT ball_on(31) AND NOT ball_on(34) AND NOT ball_on(37) AND NOT ball_on(40) AND NOT ball_on(43) AND NOT ball_on(46);
    green <= NOT ball_on(2) AND NOT ball_on(5) AND NOT ball_on(8) AND NOT ball_on(11) AND NOT cursor_on NOT ball_on(14) AND NOT ball_on(17) AND NOT ball_on(20) AND NOT ball_on(23) AND NOT ball_on(26) AND NOT ball_on(29) AND NOT ball_on(32) AND NOT ball_on(35) AND NOT ball_on(38) AND NOT ball_on(41) AND NOT ball_on(44) AND NOT ball_on(47); 

IF (pixel_col >= ballx(12) - ball_size) AND
          (pixel_col <= ballx(12) + ball_size) AND
             (pixel_row >= bally(12) - ball_size) AND
             (pixel_row <= bally(12) + ball_size) THEN
                IF (ballx(12) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(12) + ball_size >= cursor_x + cursor_size) AND
                       (bally(12) - ball_size <= cursor_y - cursor_size) AND
			           (bally(12) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(12) <= '1';END IF;
       ELSE ball_on(12) <= '0'; END IF;

IF (pixel_col >= ballx(13) - ball_size) AND
          (pixel_col <= ballx(13) + ball_size) AND
             (pixel_row >= bally(13) - ball_size) AND
             (pixel_row <= bally(13) + ball_size) THEN
                IF (ballx(13) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(13) + ball_size >= cursor_x + cursor_size) AND
                       (bally(13) - ball_size <= cursor_y - cursor_size) AND
			           (bally(13) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(13) <= '1';END IF;
       ELSE ball_on(13) <= '0'; END IF;

IF (pixel_col >= ballx(14) - ball_size) AND
          (pixel_col <= ballx(14) + ball_size) AND
             (pixel_row >= bally(14) - ball_size) AND
             (pixel_row <= bally(14) + ball_size) THEN
                IF (ballx(14) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(14) + ball_size >= cursor_x + cursor_size) AND
                       (bally(14) - ball_size <= cursor_y - cursor_size) AND
			           (bally(14) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(14) <= '1';END IF;
       ELSE ball_on(14) <= '0'; END IF;

IF (pixel_col >= ballx(15) - ball_size) AND
          (pixel_col <= ballx(15) + ball_size) AND
             (pixel_row >= bally(15) - ball_size) AND
             (pixel_row <= bally(15) + ball_size) THEN
                IF (ballx(15) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(15) + ball_size >= cursor_x + cursor_size) AND
                       (bally(15) - ball_size <= cursor_y - cursor_size) AND
			           (bally(15) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(15) <= '1';END IF;
       ELSE ball_on(15) <= '0'; END IF;

IF (pixel_col >= ballx(16) - ball_size) AND
          (pixel_col <= ballx(16) + ball_size) AND
             (pixel_row >= bally(16) - ball_size) AND
             (pixel_row <= bally(16) + ball_size) THEN
                IF (ballx(16) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(16) + ball_size >= cursor_x + cursor_size) AND
                       (bally(16) - ball_size <= cursor_y - cursor_size) AND
			           (bally(16) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(16) <= '1';END IF;
       ELSE ball_on(16) <= '0'; END IF;

IF (pixel_col >= ballx(17) - ball_size) AND
          (pixel_col <= ballx(17) + ball_size) AND
             (pixel_row >= bally(17) - ball_size) AND
             (pixel_row <= bally(17) + ball_size) THEN
                IF (ballx(17) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(17) + ball_size >= cursor_x + cursor_size) AND
                       (bally(17) - ball_size <= cursor_y - cursor_size) AND
			           (bally(17) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(17) <= '1';END IF;
       ELSE ball_on(17) <= '0'; END IF;

IF (pixel_col >= ballx(18) - ball_size) AND
          (pixel_col <= ballx(18) + ball_size) AND
             (pixel_row >= bally(18) - ball_size) AND
             (pixel_row <= bally(18) + ball_size) THEN
                IF (ballx(18) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(18) + ball_size >= cursor_x + cursor_size) AND
                       (bally(18) - ball_size <= cursor_y - cursor_size) AND
			           (bally(18) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(18) <= '1';END IF;
       ELSE ball_on(18) <= '0'; END IF;

IF (pixel_col >= ballx(19) - ball_size) AND
          (pixel_col <= ballx(19) + ball_size) AND
             (pixel_row >= bally(19) - ball_size) AND
             (pixel_row <= bally(19) + ball_size) THEN
                IF (ballx(19) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(19) + ball_size >= cursor_x + cursor_size) AND
                       (bally(19) - ball_size <= cursor_y - cursor_size) AND
			           (bally(19) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(19) <= '1';END IF;
       ELSE ball_on(19) <= '0'; END IF;

IF (pixel_col >= ballx(20) - ball_size) AND
          (pixel_col <= ballx(20) + ball_size) AND
             (pixel_row >= bally(20) - ball_size) AND
             (pixel_row <= bally(20) + ball_size) THEN
                IF (ballx(20) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(20) + ball_size >= cursor_x + cursor_size) AND
                       (bally(20) - ball_size <= cursor_y - cursor_size) AND
			           (bally(20) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(20) <= '1';END IF;
       ELSE ball_on(20) <= '0'; END IF;

IF (pixel_col >= ballx(21) - ball_size) AND
          (pixel_col <= ballx(21) + ball_size) AND
             (pixel_row >= bally(21) - ball_size) AND
             (pixel_row <= bally(21) + ball_size) THEN
                IF (ballx(21) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(21) + ball_size >= cursor_x + cursor_size) AND
                       (bally(21) - ball_size <= cursor_y - cursor_size) AND
			           (bally(21) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(21) <= '1';END IF;
       ELSE ball_on(21) <= '0'; END IF;

IF (pixel_col >= ballx(22) - ball_size) AND
          (pixel_col <= ballx(22) + ball_size) AND
             (pixel_row >= bally(22) - ball_size) AND
             (pixel_row <= bally(22) + ball_size) THEN
                IF (ballx(22) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(22) + ball_size >= cursor_x + cursor_size) AND
                       (bally(22) - ball_size <= cursor_y - cursor_size) AND
			           (bally(22) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(22) <= '1';END IF;
       ELSE ball_on(22) <= '0'; END IF;

IF (pixel_col >= ballx(23) - ball_size) AND
          (pixel_col <= ballx(23) + ball_size) AND
             (pixel_row >= bally(23) - ball_size) AND
             (pixel_row <= bally(23) + ball_size) THEN
                IF (ballx(23) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(23) + ball_size >= cursor_x + cursor_size) AND
                       (bally(23) - ball_size <= cursor_y - cursor_size) AND
			           (bally(23) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(23) <= '1';END IF;
       ELSE ball_on(23) <= '0'; END IF;

IF (pixel_col >= ballx(24) - ball_size) AND
          (pixel_col <= ballx(24) + ball_size) AND
             (pixel_row >= bally(24) - ball_size) AND
             (pixel_row <= bally(24) + ball_size) THEN
                IF (ballx(24) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(24) + ball_size >= cursor_x + cursor_size) AND
                       (bally(24) - ball_size <= cursor_y - cursor_size) AND
			           (bally(24) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(24) <= '1';END IF;
       ELSE ball_on(24) <= '0'; END IF;

IF (pixel_col >= ballx(25) - ball_size) AND
          (pixel_col <= ballx(25) + ball_size) AND
             (pixel_row >= bally(25) - ball_size) AND
             (pixel_row <= bally(25) + ball_size) THEN
                IF (ballx(25) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(25) + ball_size >= cursor_x + cursor_size) AND
                       (bally(25) - ball_size <= cursor_y - cursor_size) AND
			           (bally(25) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(25) <= '1';END IF;
       ELSE ball_on(25) <= '0'; END IF;

IF (pixel_col >= ballx(26) - ball_size) AND
          (pixel_col <= ballx(26) + ball_size) AND
             (pixel_row >= bally(26) - ball_size) AND
             (pixel_row <= bally(26) + ball_size) THEN
                IF (ballx(26) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(26) + ball_size >= cursor_x + cursor_size) AND
                       (bally(26) - ball_size <= cursor_y - cursor_size) AND
			           (bally(26) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(26) <= '1';END IF;
       ELSE ball_on(26) <= '0'; END IF;

IF (pixel_col >= ballx(27) - ball_size) AND
          (pixel_col <= ballx(27) + ball_size) AND
             (pixel_row >= bally(27) - ball_size) AND
             (pixel_row <= bally(27) + ball_size) THEN
                IF (ballx(27) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(27) + ball_size >= cursor_x + cursor_size) AND
                       (bally(27) - ball_size <= cursor_y - cursor_size) AND
			           (bally(27) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(27) <= '1';END IF;
       ELSE ball_on(27) <= '0'; END IF;

IF (pixel_col >= ballx(28) - ball_size) AND
          (pixel_col <= ballx(28) + ball_size) AND
             (pixel_row >= bally(28) - ball_size) AND
             (pixel_row <= bally(28) + ball_size) THEN
                IF (ballx(28) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(28) + ball_size >= cursor_x + cursor_size) AND
                       (bally(28) - ball_size <= cursor_y - cursor_size) AND
			           (bally(28) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(28) <= '1';END IF;
       ELSE ball_on(28) <= '0'; END IF;

IF (pixel_col >= ballx(29) - ball_size) AND
          (pixel_col <= ballx(29) + ball_size) AND
             (pixel_row >= bally(29) - ball_size) AND
             (pixel_row <= bally(29) + ball_size) THEN
                IF (ballx(29) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(29) + ball_size >= cursor_x + cursor_size) AND
                       (bally(29) - ball_size <= cursor_y - cursor_size) AND
			           (bally(29) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(29) <= '1';END IF;
       ELSE ball_on(29) <= '0'; END IF;

IF (pixel_col >= ballx(30) - ball_size) AND
          (pixel_col <= ballx(30) + ball_size) AND
             (pixel_row >= bally(30) - ball_size) AND
             (pixel_row <= bally(30) + ball_size) THEN
                IF (ballx(30) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(30) + ball_size >= cursor_x + cursor_size) AND
                       (bally(30) - ball_size <= cursor_y - cursor_size) AND
			           (bally(30) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(30) <= '1';END IF;
       ELSE ball_on(30) <= '0'; END IF;

IF (pixel_col >= ballx(31) - ball_size) AND
          (pixel_col <= ballx(31) + ball_size) AND
             (pixel_row >= bally(31) - ball_size) AND
             (pixel_row <= bally(31) + ball_size) THEN
                IF (ballx(31) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(31) + ball_size >= cursor_x + cursor_size) AND
                       (bally(31) - ball_size <= cursor_y - cursor_size) AND
			           (bally(31) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(31) <= '1';END IF;
       ELSE ball_on(31) <= '0'; END IF;

IF (pixel_col >= ballx(32) - ball_size) AND
          (pixel_col <= ballx(32) + ball_size) AND
             (pixel_row >= bally(32) - ball_size) AND
             (pixel_row <= bally(32) + ball_size) THEN
                IF (ballx(32) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(32) + ball_size >= cursor_x + cursor_size) AND
                       (bally(32) - ball_size <= cursor_y - cursor_size) AND
			           (bally(32) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(32) <= '1';END IF;
       ELSE ball_on(32) <= '0'; END IF;

IF (pixel_col >= ballx(33) - ball_size) AND
          (pixel_col <= ballx(33) + ball_size) AND
             (pixel_row >= bally(33) - ball_size) AND
             (pixel_row <= bally(33) + ball_size) THEN
                IF (ballx(33) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(33) + ball_size >= cursor_x + cursor_size) AND
                       (bally(33) - ball_size <= cursor_y - cursor_size) AND
			           (bally(33) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(33) <= '1';END IF;
       ELSE ball_on(33) <= '0'; END IF;

IF (pixel_col >= ballx(34) - ball_size) AND
          (pixel_col <= ballx(34) + ball_size) AND
             (pixel_row >= bally(34) - ball_size) AND
             (pixel_row <= bally(34) + ball_size) THEN
                IF (ballx(34) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(34) + ball_size >= cursor_x + cursor_size) AND
                       (bally(34) - ball_size <= cursor_y - cursor_size) AND
			           (bally(34) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(34) <= '1';END IF;
       ELSE ball_on(34) <= '0'; END IF;

IF (pixel_col >= ballx(35) - ball_size) AND
          (pixel_col <= ballx(35) + ball_size) AND
             (pixel_row >= bally(35) - ball_size) AND
             (pixel_row <= bally(35) + ball_size) THEN
                IF (ballx(35) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(35) + ball_size >= cursor_x + cursor_size) AND
                       (bally(35) - ball_size <= cursor_y - cursor_size) AND
			           (bally(35) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(35) <= '1';END IF;
       ELSE ball_on(35) <= '0'; END IF;

IF (pixel_col >= ballx(36) - ball_size) AND
          (pixel_col <= ballx(36) + ball_size) AND
             (pixel_row >= bally(36) - ball_size) AND
             (pixel_row <= bally(36) + ball_size) THEN
                IF (ballx(36) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(36) + ball_size >= cursor_x + cursor_size) AND
                       (bally(36) - ball_size <= cursor_y - cursor_size) AND
			           (bally(36) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(36) <= '1';END IF;
       ELSE ball_on(36) <= '0'; END IF;

IF (pixel_col >= ballx(37) - ball_size) AND
          (pixel_col <= ballx(37) + ball_size) AND
             (pixel_row >= bally(37) - ball_size) AND
             (pixel_row <= bally(37) + ball_size) THEN
                IF (ballx(37) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(37) + ball_size >= cursor_x + cursor_size) AND
                       (bally(37) - ball_size <= cursor_y - cursor_size) AND
			           (bally(37) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(37) <= '1';END IF;
       ELSE ball_on(37) <= '0'; END IF;

IF (pixel_col >= ballx(38) - ball_size) AND
          (pixel_col <= ballx(38) + ball_size) AND
             (pixel_row >= bally(38) - ball_size) AND
             (pixel_row <= bally(38) + ball_size) THEN
                IF (ballx(38) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(38) + ball_size >= cursor_x + cursor_size) AND
                       (bally(38) - ball_size <= cursor_y - cursor_size) AND
			           (bally(38) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(38) <= '1';END IF;
       ELSE ball_on(38) <= '0'; END IF;

IF (pixel_col >= ballx(39) - ball_size) AND
          (pixel_col <= ballx(39) + ball_size) AND
             (pixel_row >= bally(39) - ball_size) AND
             (pixel_row <= bally(39) + ball_size) THEN
                IF (ballx(39) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(39) + ball_size >= cursor_x + cursor_size) AND
                       (bally(39) - ball_size <= cursor_y - cursor_size) AND
			           (bally(39) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(39) <= '1';END IF;
       ELSE ball_on(39) <= '0'; END IF;

IF (pixel_col >= ballx(40) - ball_size) AND
          (pixel_col <= ballx(40) + ball_size) AND
             (pixel_row >= bally(40) - ball_size) AND
             (pixel_row <= bally(40) + ball_size) THEN
                IF (ballx(40) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(40) + ball_size >= cursor_x + cursor_size) AND
                       (bally(40) - ball_size <= cursor_y - cursor_size) AND
			           (bally(40) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(40) <= '1';END IF;
       ELSE ball_on(40) <= '0'; END IF;

IF (pixel_col >= ballx(41) - ball_size) AND
          (pixel_col <= ballx(41) + ball_size) AND
             (pixel_row >= bally(41) - ball_size) AND
             (pixel_row <= bally(41) + ball_size) THEN
                IF (ballx(41) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(41) + ball_size >= cursor_x + cursor_size) AND
                       (bally(41) - ball_size <= cursor_y - cursor_size) AND
			           (bally(41) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(41) <= '1';END IF;
       ELSE ball_on(41) <= '0'; END IF;

IF (pixel_col >= ballx(42) - ball_size) AND
          (pixel_col <= ballx(42) + ball_size) AND
             (pixel_row >= bally(42) - ball_size) AND
             (pixel_row <= bally(42) + ball_size) THEN
                IF (ballx(42) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(42) + ball_size >= cursor_x + cursor_size) AND
                       (bally(42) - ball_size <= cursor_y - cursor_size) AND
			           (bally(42) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(42) <= '1';END IF;
       ELSE ball_on(42) <= '0'; END IF;

IF (pixel_col >= ballx(43) - ball_size) AND
          (pixel_col <= ballx(43) + ball_size) AND
             (pixel_row >= bally(43) - ball_size) AND
             (pixel_row <= bally(43) + ball_size) THEN
                IF (ballx(43) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(43) + ball_size >= cursor_x + cursor_size) AND
                       (bally(43) - ball_size <= cursor_y - cursor_size) AND
			           (bally(43) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(43) <= '1';END IF;
       ELSE ball_on(43) <= '0'; END IF;

IF (pixel_col >= ballx(44) - ball_size) AND
          (pixel_col <= ballx(44) + ball_size) AND
             (pixel_row >= bally(44) - ball_size) AND
             (pixel_row <= bally(44) + ball_size) THEN
                IF (ballx(44) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(44) + ball_size >= cursor_x + cursor_size) AND
                       (bally(44) - ball_size <= cursor_y - cursor_size) AND
			           (bally(44) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(44) <= '1';END IF;
       ELSE ball_on(44) <= '0'; END IF;

IF (pixel_col >= ballx(45) - ball_size) AND
          (pixel_col <= ballx(45) + ball_size) AND
             (pixel_row >= bally(45) - ball_size) AND
             (pixel_row <= bally(45) + ball_size) THEN
                IF (ballx(45) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(45) + ball_size >= cursor_x + cursor_size) AND
                       (bally(45) - ball_size <= cursor_y - cursor_size) AND
			           (bally(45) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(45) <= '1';END IF;
       ELSE ball_on(45) <= '0'; END IF;

IF (pixel_col >= ballx(46) - ball_size) AND
          (pixel_col <= ballx(46) + ball_size) AND
             (pixel_row >= bally(46) - ball_size) AND
             (pixel_row <= bally(46) + ball_size) THEN
                IF (ballx(46) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(46) + ball_size >= cursor_x + cursor_size) AND
                       (bally(46) - ball_size <= cursor_y - cursor_size) AND
			           (bally(46) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(46) <= '1';END IF;
       ELSE ball_on(46) <= '0'; END IF;

IF (pixel_col >= ballx(47) - ball_size) AND
          (pixel_col <= ballx(47) + ball_size) AND
             (pixel_row >= bally(47) - ball_size) AND
             (pixel_row <= bally(47) + ball_size) THEN
                IF (ballx(47) - ball_size <= cursor_x - cursor_size) AND
                   (ballx(47) + ball_size >= cursor_x + cursor_size) AND
                       (bally(47) - ball_size <= cursor_y - cursor_size) AND
			           (bally(47) + ball_size >= cursor_y + cursor_size) THEN
			                ball_on(47) <= '1';END IF;
       ELSE ball_on(47) <= '0'; END IF;


